module veb

import io
import net
import net.http
import net.urllib
import os
import time
import strings
import picoev
